`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:25:09 12/08/2022 
// Design Name: 
// Module Name:    lights 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module lights(
    input a,state,next_state,a,b,c,d,
    output r1,g1,y1,r2,g2,y2,r3,g3,y3,r4,g4,y4
    );


endmodule
